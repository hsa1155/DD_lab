`include "Adder.v"
`include "BWA_add.v"
`include "BWA_EXadd.v"
module BWA(clk,a,b,ans);
	input clk;
	input [31:0]a,b;
	output [63:0] ans;
	
	wire [31:0] add0,add1,add2,add3,add4,add5,add6,add7,add8,add9,add10,add11,add12,add13,add14,add15,add16,add17,add18,add19,add20,add21,add22,add23,add24,add25,add26,add27,add28,add29,add30,add31;
	wire [63:0] abd0,abd1,abd2,abd3,abd4,abd5,abd6,abd7,abd8,abd9,abd10,abd11,abd12,abd13,abd14,abd15,abd16,abd17,abd18,abd19,abd20,abd21,abd22,abd23,abd24,abd25,abd26,abd27,abd28,abd29,abd30,abd31,abd32;
	wire [63:0] sum0,sum1,sum2,sum3,sum4,sum5,sum6,sum7,sum8,sum9,sum10,sum11,sum12,sum13,sum14,sum15,sum16,sum17,sum18,sum19,sum20,sum21,sum22,sum23,sum24,sum25,sum26,sum27,sum28,sum29,sum30,sum31;
	BWA_add Badd0(clk,a,b[0],add0);
	BWA_add Badd1(clk,a,b[1],add1);
	BWA_add Badd2(clk,a,b[2],add2);
	BWA_add Badd3(clk,a,b[3],add3);
	BWA_add Badd4(clk,a,b[4],add4);
	BWA_add Badd5(clk,a,b[5],add5);
	BWA_add Badd6(clk,a,b[6],add6);
	BWA_add Badd7(clk,a,b[7],add7);
	BWA_add Badd8(clk,a,b[8],add8);
	BWA_add Badd9(clk,a,b[9],add9);
	BWA_add Badd10(clk,a,b[10],add10);
	BWA_add Badd11(clk,a,b[11],add11);
	BWA_add Badd12(clk,a,b[12],add12);
	BWA_add Badd13(clk,a,b[13],add13);
	BWA_add Badd14(clk,a,b[14],add14);
	BWA_add Badd15(clk,a,b[15],add15);
	BWA_add Badd16(clk,a,b[16],add16);
	BWA_add Badd17(clk,a,b[17],add17);
	BWA_add Badd18(clk,a,b[18],add18);
	BWA_add Badd19(clk,a,b[19],add19);
	BWA_add Badd20(clk,a,b[20],add20);
	BWA_add Badd21(clk,a,b[21],add21);
	BWA_add Badd22(clk,a,b[22],add22);
	BWA_add Badd23(clk,a,b[23],add23);
	BWA_add Badd24(clk,a,b[24],add24);
	BWA_add Badd25(clk,a,b[25],add25);
	BWA_add Badd26(clk,a,b[26],add26);
	BWA_add Badd27(clk,a,b[27],add27);
	BWA_add Badd28(clk,a,b[28],add28);
	BWA_add Badd29(clk,a,b[29],add29);
	BWA_add Badd30(clk,a,b[30],add30);
	BWA_EXadd Badd31(clk,a,b[31],add31);
	
	assign abd0 = {32'b0, add0};
	assign abd1 = {31'b0, add1,1'b0};
	assign abd2 = {30'b0, add2,2'b0};
	assign abd3 = {29'b0, add3,3'b0};
	assign abd4 = {28'b0, add4,4'b0};
	assign abd5 = {27'b0, add5,5'b0};
	assign abd6 = {26'b0, add6,6'b0};
	assign abd7 = {25'b0, add7,7'b0};
	assign abd8 = {24'b0, add8,8'b0};
	assign abd9 = {23'b0, add9,9'b0};
	assign abd10 = {22'b0, add10,10'b0};
	assign abd11 = {21'b0, add11,11'b0};
	assign abd12 = {20'b0, add12,12'b0};
	assign abd13 = {19'b0, add13,13'b0};
	assign abd14 = {18'b0, add14,14'b0};
	assign abd15 = {17'b0, add15,15'b0};
	assign abd16 = {16'b0, add16,16'b0};
	assign abd17 = {15'b0, add17,17'b0};
	assign abd18 = {14'b0, add18,18'b0};
	assign abd19 = {13'b0, add19,19'b0};
	assign abd20 = {12'b0, add20,20'b0};
	assign abd21 = {11'b0, add21,21'b0};
	assign abd22 = {10'b0, add22,22'b0};
	assign abd23 = {9'b0, add23,23'b0};
	assign abd24 = {8'b0, add24,24'b0};
	assign abd25 = {7'b0, add25,25'b0};
	assign abd26 = {6'b0, add26,26'b0};
	assign abd27 = {5'b0, add27,27'b0};
	assign abd28 = {4'b0, add28,28'b0};
	assign abd29 = {3'b0, add29,29'b0};
	assign abd30 = {2'b0, add30,30'b0};
	assign abd31 = {1'b0, add31,31'b0};
	assign abd32 = {1'b1,30'b0,1'b1,32'b0};
	adder adder1(clk,abd0,abd1,sum0);
	adder adder2(clk,sum0,abd2,sum1);
	adder adder3(clk,sum1,abd3,sum2);
	adder adder4(clk,sum2,abd4,sum3);
	adder adder5(clk,sum3,abd5,sum4);
	adder adder6(clk,sum4,abd6,sum5);
	adder adder7(clk,sum5,abd7,sum6);
	adder adder8(clk,sum6,abd8,sum7);
	adder adder9(clk,sum7,abd9,sum8);
	adder adder10(clk,sum8,abd10,sum9);
	adder adder11(clk,sum9,abd11,sum10);
	adder adder12(clk,sum10,abd12,sum11);
	adder adder13(clk,sum11,abd13,sum12);
	adder adder14(clk,sum12,abd14,sum13);
	adder adder15(clk,sum13,abd15,sum14);
	adder adder16(clk,sum14,abd16,sum15);
	adder adder17(clk,sum15,abd17,sum16);
	adder adder18(clk,sum16,abd18,sum17);
	adder adder19(clk,sum17,abd19,sum18);
	adder adder20(clk,sum18,abd20,sum19);
	adder adder21(clk,sum19,abd21,sum20);
	adder adder22(clk,sum20,abd22,sum21);
	adder adder23(clk,sum21,abd23,sum22);
	adder adder24(clk,sum22,abd24,sum23);
	adder adder25(clk,sum23,abd25,sum24);
	adder adder26(clk,sum24,abd26,sum25);
	adder adder27(clk,sum25,abd27,sum26);
	adder adder28(clk,sum26,abd28,sum27);
	adder adder29(clk,sum27,abd29,sum28);
	adder adder30(clk,sum28,abd30,sum29);
	adder adder31(clk,sum29,abd31,sum30);
	adder adder32(clk,sum30,abd32,ans);
endmodule
