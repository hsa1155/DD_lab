module BWA_add(clk,a,b,out);
	input clk;
	input [31:0] a;
	input b;
	output [31:0] out;
	assign out[0] = a[0]&b;
	assign out[1] = a[1]&b;
	assign out[2] = a[2]&b;
	assign out[3] = a[3]&b;
	assign out[4] = a[4]&b;
	assign out[5] = a[5]&b;
	assign out[6] = a[6]&b;
	assign out[7] = a[7]&b;
	assign out[8] = a[8]&b;
	assign out[9] = a[9]&b;
	assign out[10] = a[10]&b;
	assign out[11] = a[11]&b;
	assign out[12] = a[12]&b;
	assign out[13] = a[13]&b;
	assign out[14] = a[14]&b;
	assign out[15] = a[15]&b;
	assign out[16] = a[16]&b;
	assign out[17] = a[17]&b;
	assign out[18] = a[18]&b;
	assign out[19] = a[19]&b;
	assign out[20] = a[20]&b;
	assign out[21] = a[21]&b;
	assign out[22] = a[22]&b;
	assign out[23] = a[23]&b;
	assign out[24] = a[24]&b;
	assign out[25] = a[25]&b;
	assign out[26] = a[26]&b;
	assign out[27] = a[27]&b;
	assign out[28] = a[28]&b;
	assign out[29] = a[29]&b;
	assign out[30] = a[30]&b;
	assign out[31] = !(a[31]&b);

endmodule